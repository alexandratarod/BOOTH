module xor_m_c3( 
  input m, c3,
  output out);
  
  
  assign out = m ^ c3;

endmodule

